//  ------------------------------------------------------------------------
// File :                       sem_task.v
// Author :                     superboy
// Created date :               2022/09/10
// Abstract     :               Unique module for record and tell the core what to do next. It will be designed upon the specific application scenarios.
// Last modified date :         2022/09/10
// -------------------------------------------------------------------
// -------------------------------------------------------------------